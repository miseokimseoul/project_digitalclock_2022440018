`timescale 1us/1us

module tb_TimerController;

    // DUT �Է�
    reg clk_1k;
    reg tick_1hz;
    reg timer_sw;

    reg btn_h_inc;
    reg btn_m_inc;
    reg btn_s_inc;
    reg btn_confirm;
    reg btn_start;
    reg btn_clear;
    reg btn_add5;
    reg btn_add10;
    reg btn_add15;

    // DUT ���
    wire [3:0] tm_h_tens;
    wire [3:0] tm_h_ones;
    wire [3:0] tm_m_tens;
    wire [3:0] tm_m_ones;
    wire [3:0] tm_s_tens;
    wire [3:0] tm_s_ones;

    wire [1:0] timer_state;
    wire       led_1_blink;
    wire [2:0] rgb_pwm;
    wire       piezo_out;
    wire [3:0] sand_count;

    // DUT �ν��Ͻ�
    TimerController dut (
        .clk_1k      (clk_1k),
        .tick_1hz    (tick_1hz),
        .timer_sw    (timer_sw),
        .btn_h_inc   (btn_h_inc),
        .btn_m_inc   (btn_m_inc),
        .btn_s_inc   (btn_s_inc),
        .btn_confirm (btn_confirm),
        .btn_start   (btn_start),
        .btn_clear   (btn_clear),
        .btn_add5    (btn_add5),
        .btn_add10   (btn_add10),
        .btn_add15   (btn_add15),
        .tm_h_tens   (tm_h_tens),
        .tm_h_ones   (tm_h_ones),
        .tm_m_tens   (tm_m_tens),
        .tm_m_ones   (tm_m_ones),
        .tm_s_tens   (tm_s_tens),
        .tm_s_ones   (tm_s_ones),
        .timer_state (timer_state),
        .led_1_blink (led_1_blink),
        .rgb_pwm     (rgb_pwm),
        .piezo_out   (piezo_out),
        .sand_count  (sand_count)
    );

    //--------------------------------------------------
    // 1 kHz Ŭ��
    //--------------------------------------------------
    initial clk_1k = 0;
    always #500 clk_1k = ~clk_1k;  // 1kHz

    //--------------------------------------------------
    // 1 Hz tick
    //--------------------------------------------------
    task tick_once;
    begin
        tick_1hz = 1'b1;
        @(posedge clk_1k);
        tick_1hz = 1'b0;
        @(posedge clk_1k);
    end
    endtask

    task tick_many;
        input integer n;
        integer i;
    begin
        for (i = 0; i < n; i = i + 1)
            tick_once();
    end
    endtask

    //--------------------------------------------------
    // ��ư �ʱ�ȭ & ���� ��ư task
    //--------------------------------------------------
    task clear_buttons;
    begin
        btn_h_inc   = 0;
        btn_m_inc   = 0;
        btn_s_inc   = 0;
        btn_confirm = 0;
        btn_start   = 0;
        btn_clear   = 0;
        btn_add5    = 0;
        btn_add10   = 0;
        btn_add15   = 0;
    end
    endtask

    task press_s_inc;
    begin
        btn_s_inc = 1;
        @(posedge clk_1k);
        btn_s_inc = 0;
        @(posedge clk_1k);
    end
    endtask

    task press_start;
    begin
        btn_start = 1;
        @(posedge clk_1k);
        btn_start = 0;
        @(posedge clk_1k);
    end
    endtask

    //--------------------------------------------------
    // ���� �ùķ��̼�
    //--------------------------------------------------
    initial begin
        tick_1hz = 0;
        timer_sw = 0;
        clear_buttons();

        // -------------------------------
        // �� ���� �ʱ�ȭ : btn_clear �޽�
        // -------------------------------
        // �ùķ��̼� ���� ���� �� Ŭ�� ���� clear=1�� ����
        // timer_state, cnt_hour/min/sec ���� 0���� ���� �ʱ�ȭ
        btn_clear = 1;
        repeat(5) @(posedge clk_1k);
        btn_clear = 0;
        repeat(5) @(posedge clk_1k);

        //--------------------------------------------------
        // [���� 1] 5�� Ÿ�̸� �� ī��Ʈ�ٿ� �� RINGING
        //--------------------------------------------------
        timer_sw = 1;
        repeat(5) @(posedge clk_1k);

        // 00:00:05 ����
        repeat(5) press_s_inc();   // tm_s = 05

        // START
        press_start();
        repeat(5) @(posedge clk_1k);

        // 5 �� 0 ī��Ʈ�ٿ� + RINGING ����
        tick_many(6);  // S_RUNNING �� S_RINGING

        // ���� ���� 3�� (piezo_out ��� Ȯ��)
        tick_many(3);

        #5000;  // ���� ����

        //--------------------------------------------------
        // [���� 2] 20�� Ÿ�̸� �� ��׶��� ����
        //--------------------------------------------------
        // �ٽ� �ѹ� clear�� �ʱ�ȭ
        btn_clear = 1;
        repeat(5) @(posedge clk_1k);
        btn_clear = 0;
        repeat(5) @(posedge clk_1k);

        timer_sw = 1;
        repeat(5) @(posedge clk_1k);

        // 00:00:20 ����
        repeat(20) press_s_inc();

        // START
        press_start();
        repeat(5) @(posedge clk_1k);

        // Ÿ�̸� ��忡�� 2�� ī��Ʈ�ٿ�
        tick_many(2);  // 20 �� 18��

        // timer_sw=0���� ���� �⺻ �ð� ��� ���� (��׶��� ����)
        timer_sw = 0;

        // ���� 18�� ���� ī��Ʈ�ٿ� �� sand_count, rgb_pwm, led_1_blink Ȯ��
        tick_many(18);

        #5000;
        $stop;
    end

endmodule
